module div2 (A, B, C, D, Out);
	input A, B, C, D;
	output Out;
	
	not inv1(Out,D);
endmodule
